package cea861d_1080p30_pkg;

parameter int TOTAL_X                     = 2200;
parameter int TOTAL_Y                     = 1125;
parameter int DE_NEGEDGE_TO_HSYNC_POSEDGE = 88;
parameter int HSYNC_WIDTH                 = 44;
parameter int HSYNC_NEGEDGE_TO_DE_POSEDGE = 148;
parameter int ACTIVE_X                    = 1920;
parameter int VERTICAL_BLNAKING_PRE       = 41;
parameter int VERTICAL_BLANKING_POST      = 4;
parameter int ACTIVE_LINES                = 1080;
parameter int VSYNC_WIDTH                 = 5;

endpackage
